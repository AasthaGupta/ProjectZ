package neuron_types is
	type neuron_in is array(8 downto 0) of bit_vector(39 downto 0);
end package;