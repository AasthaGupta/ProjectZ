package neuron_types is
	type network_vector is array(0 to 8) of bit_vector(39 downto 0);
end package;
